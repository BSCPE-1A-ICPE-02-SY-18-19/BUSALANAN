CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 108 189 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6295 0 0
2
43530.5 0
0
9 CC 7-Seg~
183 842 166 0 18 19
10 12 11 10 5 4 3 2 18 19
0 0 0 1 1 1 1 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
332 0 0
2
43530.5 1
0
9 2-In AND~
219 545 49 0 3 22
0 14 7 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9737 0 0
2
43530.5 2
0
9 2-In AND~
219 390 52 0 3 22
0 9 8 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9910 0 0
2
43530.5 3
0
6 74112~
219 604 225 0 7 32
0 17 13 15 13 17 20 6
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3834 0 0
2
43530.5 4
0
6 74112~
219 504 226 0 7 32
0 17 14 15 14 17 21 7
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3138 0 0
2
43530.5 5
0
6 74112~
219 395 231 0 7 32
0 17 9 15 9 17 22 8
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
5409 0 0
2
43530.5 6
0
6 74112~
219 289 231 0 7 32
0 17 16 15 16 17 23 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
983 0 0
2
43530.5 7
0
6 74LS48
188 761 246 0 14 29
0 6 7 8 9 24 25 2 3 4
5 10 11 12 26
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6652 0 0
2
43530.5 8
0
2 +V
167 131 125 0 1 3
0 17
0
0 0 54256 0
2 5V
-6 -22 8 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4281 0 0
2
43530.5 9
0
7 Pulser~
4 70 313 0 10 12
0 27 28 15 29 0 0 5 5 5
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6847 0 0
2
43530.5 10
0
35
7 7 2 0 0 4224 0 9 2 0 0 3
793 210
857 210
857 202
8 6 3 0 0 4224 0 9 2 0 0 3
793 219
851 219
851 202
9 5 4 0 0 4224 0 9 2 0 0 3
793 228
845 228
845 202
10 4 5 0 0 4224 0 9 2 0 0 3
793 237
839 237
839 202
7 1 6 0 0 12416 0 5 9 0 0 4
628 189
675 189
675 210
729 210
2 0 7 0 0 12416 0 9 0 0 14 5
729 219
705 219
705 116
530 116
530 159
0 3 8 0 0 8320 0 0 9 18 0 5
425 248
425 323
717 323
717 228
729 228
0 7 9 0 0 4096 0 0 8 24 0 2
329 195
313 195
11 3 10 0 0 8320 0 9 2 0 0 3
793 246
833 246
833 202
12 2 11 0 0 8320 0 9 2 0 0 3
793 255
827 255
827 202
13 1 12 0 0 8320 0 9 2 0 0 3
793 264
821 264
821 202
0 4 13 0 0 4096 0 0 5 13 0 3
566 95
566 207
580 207
3 2 13 0 0 8320 0 3 5 0 0 3
566 49
566 189
580 189
2 7 7 0 0 0 0 3 6 0 0 6
521 58
512 58
512 159
539 159
539 190
528 190
0 4 14 0 0 4224 0 0 6 17 0 3
429 52
429 208
480 208
0 1 14 0 0 0 0 0 3 17 0 3
465 52
465 40
521 40
3 2 14 0 0 0 0 4 6 0 0 4
411 52
466 52
466 190
480 190
2 7 8 0 0 0 0 4 7 0 0 6
366 61
356 61
356 248
433 248
433 195
419 195
1 0 9 0 0 8192 0 4 0 0 24 3
366 43
335 43
335 195
3 0 15 0 0 8192 0 5 0 0 21 4
574 198
570 198
570 304
470 304
3 0 15 0 0 12288 0 6 0 0 22 4
474 199
470 199
470 304
361 304
3 0 15 0 0 12288 0 7 0 0 25 4
365 204
361 204
361 304
251 304
0 4 9 0 0 0 0 0 7 24 0 3
343 195
343 213
371 213
4 2 9 0 0 12416 0 9 7 0 0 6
729 237
705 237
705 286
326 286
326 195
371 195
3 3 15 0 0 4224 0 11 8 0 0 4
94 304
251 304
251 204
259 204
0 4 16 0 0 8192 0 0 8 27 0 3
144 189
144 213
265 213
1 2 16 0 0 4224 0 1 8 0 0 4
120 189
251 189
251 195
265 195
5 0 17 0 0 8192 0 8 0 0 31 3
289 243
289 272
395 272
5 0 17 0 0 12288 0 5 0 0 32 5
604 237
604 272
648 272
648 136
604 136
5 0 17 0 0 0 0 6 0 0 29 3
504 238
504 272
604 272
5 0 17 0 0 0 0 7 0 0 30 3
395 243
395 272
504 272
0 1 17 0 0 0 0 0 5 33 0 3
504 136
604 136
604 162
0 1 17 0 0 0 0 0 6 34 0 3
395 136
504 136
504 163
1 0 17 0 0 0 0 7 0 0 35 3
395 168
395 134
289 134
1 1 17 0 0 4224 0 10 8 0 0 3
131 134
289 134
289 168
1
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 21
168 354 325 381
180 362 312 381
21 Busalanan, Harold Gil
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
